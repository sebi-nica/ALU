module div_logic(
    input[3:0] state_curr,
    input cnt_done, q0, a7,
    output[3:0] state_nxt,
    output c0, c1, c2, c3, c4, c5, c6, c7
);

    assign state_curr[0] =
    assign state_curr[1] =
    assign state_curr[2] =
    assign state_curr[3] =
    assign c0 =
    assign c1 =
    assign c2 =
    assign c3 =
    assign c4 =
    assign c5 =
    assign c6 =
    assign c7 =
endmodule